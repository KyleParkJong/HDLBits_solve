module top_module (
    input [99:0] a, b, 
    input cin,
    output [99:0] cout, sum
);
    

endmodule
